library ieee;
use ieee.std_logic_1164.all;

entity phelmino_core is
  
  port (
    -- Clock and reset signals
    clk	  : in std_logic;
    rst_n : in std_logic);

end entity phelmino_core;
